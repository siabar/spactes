20059004|_SUG_Arteria_afectada|a. basilar|Arteria basilar|no
20059004|_SUG_Arteria_afectada|a.basilar|Arteria basilar|si
20059004|_SUG_Arteria_afectada|ab|Arteria basilar|no
20059004|_SUG_Arteria_afectada|art basilar|Arteria basilar|no
20059004|_SUG_Arteria_afectada|arteria basilar|Arteria basilar|no
20059004|_SUG_Arteria_afectada|acc|Arteria carótida común|no
20059004|_SUG_Arteria_afectada|arteria acc|Arteria carótida común|no
20059004|_SUG_Arteria_afectada|arteria carotida comun|Arteria carótida común|no
20059004|_SUG_Arteria_afectada|carotide|Arteria carótida común|no
20059004|_SUG_Arteria_afectada|arteria carotide|Arteria carótida común|no
20059004|_SUG_Arteria_afectada|arteria carotidea|Arteria carótida común|no
20059004|_SUG_Arteria_afectada|arteria carotidi|Arteria carótida común|no
20059004|_SUG_Arteria_afectada|carotida|Arteria carótida común|no
20059004|_SUG_Arteria_afectada|a. carotida interna|Arteria carótida interna|no
20059004|_SUG_Arteria_afectada|a.carotida interna|Arteria carótida interna|no
20059004|_SUG_Arteria_afectada|aci|Arteria carótida interna|no
20059004|_SUG_Arteria_afectada|arteria aci|Arteria carótida interna|no
20059004|_SUG_Arteria_afectada|arteria carotida interna|Arteria carótida interna|no
20059004|_SUG_Arteria_afectada|arteria ica|Arteria carótida interna|no
20059004|_SUG_Arteria_afectada|carotida interna|Arteria carótida interna|no
20059004|_SUG_Arteria_afectada|ica|Arteria carótida interna|no
20059004|_SUG_Arteria_afectada|arteria c1|Arteria carótida interna segmento cervical o C1|no
20059004|_SUG_Arteria_afectada|c1|Arteria carótida interna segmento cervical o C1|no
20059004|_SUG_Arteria_afectada|aci-t|Arteria carótida interna terminal (o ACI-T/ TICA)|no
20059004|_SUG_Arteria_afectada|arteria aci-t|Arteria carótida interna terminal (o ACI-T/ TICA)|no
20059004|_SUG_Arteria_afectada|arteria carotida interna terminal|Arteria carótida interna terminal (o ACI-T/ TICA)|no
20059004|_SUG_Arteria_afectada|arteria tica|Arteria carótida interna terminal (o ACI-T/ TICA)|no
20059004|_SUG_Arteria_afectada|tica|Arteria carótida interna terminal (o ACI-T/ TICA)|no
20059004|_SUG_Arteria_afectada|arteria carotida primitiva|Arteria carótida primitiva|no
20059004|_SUG_Arteria_afectada|carotida primitiva|Arteria carótida primitiva|no
20059004|_SUG_Arteria_afectada|aica|Arteria cerebelosa posteroinferior (o PICA)|no
20059004|_SUG_Arteria_afectada|arteria aica|Arteria cerebelosa posteroinferior (o PICA)|no
20059004|_SUG_Arteria_afectada|arteria cerebelosa anteroinferior|Arteria cerebelosa posteroinferior (o PICA)|no
20059004|_SUG_Arteria_afectada|arteria cerebelosa posteroinferior|Arteria cerebelosa posteroinferior (o PICA)|no
20059004|_SUG_Arteria_afectada|arteria cerebelosa superior|Arteria cerebelosa posteroinferior (o PICA)|no
20059004|_SUG_Arteria_afectada|arteria pica|Arteria cerebelosa posteroinferior (o PICA)|no
20059004|_SUG_Arteria_afectada|pica|Arteria cerebelosa posteroinferior (o PICA)|no
20059004|_SUG_Arteria_afectada|acs|Arteria cerebelosa superior|no
20059004|_SUG_Arteria_afectada|arteria acs|Arteria cerebelosa superior|no
20059004|_SUG_Arteria_afectada|aca|Arteria cerebral anterior|no
20059004|_SUG_Arteria_afectada|acoa|Arteria cerebral anterior|no
20059004|_SUG_Arteria_afectada|arteria aca|Arteria cerebral anterior|no
20059004|_SUG_Arteria_afectada|arteria acoa|Arteria cerebral anterior|no
20059004|_SUG_Arteria_afectada|arteria cerebral anterior|Arteria cerebral anterior|no
20059004|_SUG_Arteria_afectada|a2|Arteria cerebral anterior segmento A2|no
20059004|_SUG_Arteria_afectada|arteria a2|Arteria cerebral anterior segmento A2|no
20059004|_SUG_Arteria_afectada|acm|Arteria cerebral media|no
20059004|_SUG_Arteria_afectada|art cerebral media|Arteria cerebral media|no
20059004|_SUG_Arteria_afectada|art. cerebral media|Arteria cerebral media|no
20059004|_SUG_Arteria_afectada|arteria acm|Arteria cerebral media|no
20059004|_SUG_Arteria_afectada|arteria cerebral media|Arteria cerebral media|no
20059004|_SUG_Arteria_afectada|arteria cerebral mitja|Arteria cerebral media|no
20059004|_SUG_Arteria_afectada|arteria cerebrals mitges|Arteria cerebral media|no
20059004|_SUG_Arteria_afectada|arteria nucleo lenticular|Arteria cerebral media|no
20059004|_SUG_Arteria_afectada|nucleo lenticular|Arteria cerebral media|no
20059004|_SUG_Arteria_afectada|arteria cerebral media segmento|Arteria cerebral media segmento|no
20059004|_SUG_Arteria_afectada|arteria m1|Arteria cerebral media segmento M1|no
20059004|_SUG_Arteria_afectada|m1|Arteria cerebral media segmento M1|no
20059004|_SUG_Arteria_afectada|arteria m2|Arteria cerebral media segmento M2|no
20059004|_SUG_Arteria_afectada|m2|Arteria cerebral media segmento M2|no
20059004|_SUG_Arteria_afectada|arteria m3|Arteria cerebral media segmento M3|no
20059004|_SUG_Arteria_afectada|m3|Arteria cerebral media segmento M3|no
20059004|_SUG_Arteria_afectada|arteria m4|Arteria cerebral media segmento M4|no
20059004|_SUG_Arteria_afectada|m4|Arteria cerebral media segmento M4|no
20059004|_SUG_Arteria_afectada|arteria m5|Arteria cerebral media segmento M5|no
20059004|_SUG_Arteria_afectada|m5|Arteria cerebral media segmento M5|no
20059004|_SUG_Arteria_afectada|arteria m6|Arteria cerebral media segmento M6|no
20059004|_SUG_Arteria_afectada|m6|Arteria cerebral media segmento M6|no
20059004|_SUG_Arteria_afectada|acp|Arteria cerebral posterior|no
20059004|_SUG_Arteria_afectada|arteria acp|Arteria cerebral posterior|no
20059004|_SUG_Arteria_afectada|arteria cerebral posterior|Arteria cerebral posterior|no
20059004|_SUG_Arteria_afectada|arteria cerebrales posteriores|Arteria cerebral posterior|no
20059004|_SUG_Arteria_afectada|cerebrales posteriores|Arteria cerebral posterior|no
20059004|_SUG_Arteria_afectada|a. circunferencial corta|Arteria circunferencial corta|no
20059004|_SUG_Arteria_afectada|a.circunferencial corta|Arteria circunferencial corta|no
20059004|_SUG_Arteria_afectada|a. coroidea ant|Arteria coroidea anterior|no
20059004|_SUG_Arteria_afectada|a.coroidea ant|Arteria coroidea anterior|no
20059004|_SUG_Arteria_afectada|arteria coroidea anterior|Arteria coroidea anterior|no
20059004|_SUG_Arteria_afectada|arteria coroidea posterior|Arteria coroidea posterior|no
20059004|_SUG_Arteria_afectada|arteria lenticular estriadas|Arteria lenticuloestriada|no
20059004|_SUG_Arteria_afectada|arteria lenticular-estriadas|Arteria lenticuloestriada|no
20059004|_SUG_Arteria_afectada|arteria lenticuloestriada|Arteria lenticuloestriada|no
20059004|_SUG_Arteria_afectada|lenticular estriadas|Arteria lenticuloestriada|no
20059004|_SUG_Arteria_afectada|lenticular-estriadas|Arteria lenticuloestriada|no
20059004|_SUG_Arteria_afectada|a. paramedia|Arteria paramedia|no
20059004|_SUG_Arteria_afectada|art. paramedia|Arteria paramedia|no
20059004|_SUG_Arteria_afectada|arteria paramedia|Arteria paramedia|no
20059004|_SUG_Arteria_afectada|arteria paramediana|Arteria paramediana|no
20059004|_SUG_Arteria_afectada|art vertebral|Arteria vertebral|no
20059004|_SUG_Arteria_afectada|arteria vertebral|Arteria vertebral|no
20059004|_SUG_Arteria_afectada|arteria v1|Arteria vertebral segmento V1|no
20059004|_SUG_Arteria_afectada|v1|Arteria vertebral segmento V1|no
20059004|_SUG_Arteria_afectada|arteria indeterm i na do|Indeterminado|no
20059004|_SUG_Arteria_afectada|arteria indeterminado|Indeterminado|no
20059004|_SUG_Arteria_afectada|arteria no especif.|Indeterminado|no
20059004|_SUG_Arteria_afectada|arteria territorio indeterminado|Indeterminado|no
20059004|_SUG_Arteria_afectada|indeterm i na do|Indeterminado|no
20059004|_SUG_Arteria_afectada|indeterminado|Indeterminado|no
20059004|_SUG_Arteria_afectada|no especif.|Indeterminado|no
20059004|_SUG_Arteria_afectada|territorio indeterminado|Indeterminado|no
20059004|_SUG_Arteria_afectada|arteria vb|Sistema vértebrobasilar|no
20059004|_SUG_Arteria_afectada|arteria vertebr basilar|Sistema vértebrobasilar|no
20059004|_SUG_Arteria_afectada|arteria vertebro basilar|Sistema vértebrobasilar|no
20059004|_SUG_Arteria_afectada|arteria vertebro-basilar|Sistema vértebrobasilar|no
20059004|_SUG_Arteria_afectada|vertebro basilar|Sistema vértebrobasilar|no
20059004|_SUG_Arteria_afectada|arteria vertebrobasilar|Sistema vértebrobasilar|no
20059004|_SUG_Arteria_afectada|vb|Sistema vértebrobasilar|no
00000010|_SUG_ASPECTS|aspects 0|ASPECTS|no
00000010|_SUG_ASPECTS|aspects score 0|ASPECTS|no
266257000|_SUG_Ataque_isquemico_transitorio|accidente transitori isquemia|Ataque isquémico transitorio|no
266257000|_SUG_Ataque_isquemico_transitorio|ait|Ataque isquémico transitorio|no
266257000|_SUG_Ataque_isquemico_transitorio|aits|Ataque isquémico transitorio|no
266257000|_SUG_Ataque_isquemico_transitorio|ataque isquemia transitorio|Ataque isquémico transitorio|no
266257000|_SUG_Ataque_isquemico_transitorio|ictus isquemia minor|Ataque isquémico transitorio|no
266257000|_SUG_Ataque_isquemico_transitorio|ictus minor|Ataque isquémico transitorio|no
266257000|_SUG_Ataque_isquemico_transitorio|infarto clinicamente regresivo|Ataque isquémico transitorio|no
266257000|_SUG_Ataque_isquemico_transitorio|isquemia cerebral transitoria|Ataque isquémico transitorio|no
266257000|_SUG_Ataque_isquemico_transitorio|tia|Ataque isquémico transitorio|no
134198009|_SUG_Etiologia|aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|causa aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|causa posiblemente aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|causa probablemente aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|de origen aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|de origen posiblemente aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|de origen probablemente aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|etiologia aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|etiologia posiblemente aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|etiologia probablemente aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|origen aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|origen posiblemente aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|origen probablemente aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|perfil aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|perfil posiblemente aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|perfil probablemente aneurisma|Aneurisma|no
134198009|_SUG_Etiologia|angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|causa angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|causa angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|causa posiblemente angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|causa posiblemente angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|causa probablemente angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|causa probablemente angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|de origen angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|de origen angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|de origen posiblemente angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|de origen posiblemente angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|de origen probablemente angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|de origen probablemente angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|etiologia angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|etiologia angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|etiologia posiblemente angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|etiologia posiblemente angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|etiologia probablemente angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|etiologia probablemente angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|origen angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|origen angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|origen posiblemente angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|origen posiblemente angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|origen probablemente angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|origen probablemente angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|perfil angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|perfil angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|perfil posiblemente angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|perfil posiblemente angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|perfil probablemente angiopatia amiloide|Angiopatía amiloide|no
134198009|_SUG_Etiologia|perfil probablemente angiopatia amiloide cerebral|Angiopatía amiloide|no
134198009|_SUG_Etiologia|ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|causa ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|causa aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|causa aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|causa posiblemente ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|causa posiblemente aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|causa posiblemente aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|causa probablemente ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|causa probablemente aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|causa probablemente aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|de origen ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|de origen aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|de origen aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|de origen posiblemente ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|de origen posiblemente aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|de origen posiblemente aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|de origen probablemente ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|de origen probablemente aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|de origen probablemente aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|etiologia ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|etiologia aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|etiologia aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|etiologia posiblemente ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|etiologia posiblemente aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|etiologia posiblemente aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|etiologia probablemente ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|etiologia probablemente aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|etiologia probablemente aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|origen ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|origen aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|origen aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|origen posiblemente ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|origen posiblemente aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|origen posiblemente aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|origen probablemente ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|origen probablemente aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|origen probablemente aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|perfil ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|perfil aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|perfil aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|perfil posiblemente ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|perfil posiblemente aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|perfil posiblemente aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|perfil probablemente ateromatosis|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|perfil probablemente aterosclerotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|perfil probablemente aterotrombotico|Aterotrombótico/aterosclerótico|no
134198009|_SUG_Etiologia|cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa embolica|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa posiblemente cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa posiblemente cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa posiblemente cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa posiblemente ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa posiblemente embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa posiblemente embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa posiblemente mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa probablemente cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa probablemente cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa probablemente cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa probablemente ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa probablemente embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa probablemente embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa probablemente mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen posiblemente cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen posiblemente cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen posiblemente cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen posiblemente ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen posiblemente embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen posiblemente embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen posiblemente mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen probablemente cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen probablemente cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen probablemente cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen probablemente ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen probablemente embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen probablemente embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|de origen probablemente mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|embolica|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia posiblemente cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia posiblemente cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia posiblemente cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia posiblemente ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia posiblemente embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia posiblemente embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia posiblemente mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia probablemente cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia probablemente cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia probablemente cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia probablemente ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia probablemente embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia probablemente embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|etiologia probablemente mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen posiblemente cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen posiblemente cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen posiblemente cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen posiblemente ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen posiblemente embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen posiblemente embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen posiblemente mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen probablemente cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen probablemente cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen probablemente cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen probablemente ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen probablemente embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen probablemente embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|origen probablemente mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil posiblemente cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil posiblemente cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil posiblemente cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil posiblemente ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil posiblemente embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil posiblemente embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil posiblemente mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil probablemente cardiaco|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil probablemente cardio embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil probablemente cardioemebolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil probablemente ce|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil probablemente embolico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil probablemente embolismo paradojico|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|perfil probablemente mecanisme embolic|Cardioembólico (CE)|no
134198009|_SUG_Etiologia|causa hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|causa posiblemente hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|causa probablemente hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|de origen hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|de origen posiblemente hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|de origen probablemente hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|etiologia hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|etiologia posiblemente hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|etiologia probablemente hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|origen hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|origen posiblemente hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|origen probablemente hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|perfil hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|perfil posiblemente hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|perfil probablemente hipertensivo|Hipertensiva|no
134198009|_SUG_Etiologia|a estudio|Indeterminada|no
134198009|_SUG_Etiologia|causa a estudio|Indeterminada|no
134198009|_SUG_Etiologia|causa no determinada|Indeterminada|no
134198009|_SUG_Etiologia|causa por determinar|Indeterminada|no
134198009|_SUG_Etiologia|causa posiblemente a estudio|Indeterminada|no
134198009|_SUG_Etiologia|causa posiblemente no determinada|Indeterminada|no
134198009|_SUG_Etiologia|causa posiblemente por determinar|Indeterminada|no
134198009|_SUG_Etiologia|causa probablemente a estudio|Indeterminada|no
134198009|_SUG_Etiologia|causa probablemente no determinada|Indeterminada|no
134198009|_SUG_Etiologia|causa probablemente por determinar|Indeterminada|no
134198009|_SUG_Etiologia|de origen a estudio|Indeterminada|no
134198009|_SUG_Etiologia|de origen no determinada|Indeterminada|no
134198009|_SUG_Etiologia|de origen por determinar|Indeterminada|no
134198009|_SUG_Etiologia|de origen posiblemente a estudio|Indeterminada|no
134198009|_SUG_Etiologia|de origen posiblemente no determinada|Indeterminada|no
134198009|_SUG_Etiologia|de origen posiblemente por determinar|Indeterminada|no
134198009|_SUG_Etiologia|de origen probablemente a estudio|Indeterminada|no
134198009|_SUG_Etiologia|de origen probablemente no determinada|Indeterminada|no
134198009|_SUG_Etiologia|de origen probablemente por determinar|Indeterminada|no
134198009|_SUG_Etiologia|etiologia a estudio|Indeterminada|no
134198009|_SUG_Etiologia|etiologia no determinada|Indeterminada|no
134198009|_SUG_Etiologia|etiologia por determinar|Indeterminada|no
134198009|_SUG_Etiologia|etiologia posiblemente a estudio|Indeterminada|no
134198009|_SUG_Etiologia|etiologia posiblemente no determinada|Indeterminada|no
134198009|_SUG_Etiologia|etiologia posiblemente por determinar|Indeterminada|no
134198009|_SUG_Etiologia|etiologia probablemente a estudio|Indeterminada|no
134198009|_SUG_Etiologia|etiologia probablemente no determinada|Indeterminada|no
134198009|_SUG_Etiologia|etiologia probablemente por determinar|Indeterminada|no
134198009|_SUG_Etiologia|no determinada|Indeterminada|no
134198009|_SUG_Etiologia|origen a estudio|Indeterminada|no
134198009|_SUG_Etiologia|origen no determinada|Indeterminada|no
134198009|_SUG_Etiologia|origen por determinar|Indeterminada|no
134198009|_SUG_Etiologia|origen posiblemente a estudio|Indeterminada|no
134198009|_SUG_Etiologia|origen posiblemente no determinada|Indeterminada|no
134198009|_SUG_Etiologia|origen posiblemente por determinar|Indeterminada|no
134198009|_SUG_Etiologia|origen probablemente a estudio|Indeterminada|no
134198009|_SUG_Etiologia|origen probablemente no determinada|Indeterminada|no
134198009|_SUG_Etiologia|origen probablemente por determinar|Indeterminada|no
134198009|_SUG_Etiologia|perfil a estudio|Indeterminada|no
134198009|_SUG_Etiologia|perfil no determinada|Indeterminada|no
134198009|_SUG_Etiologia|perfil por determinar|Indeterminada|no
134198009|_SUG_Etiologia|perfil posiblemente a estudio|Indeterminada|no
134198009|_SUG_Etiologia|perfil posiblemente no determinada|Indeterminada|no
134198009|_SUG_Etiologia|perfil posiblemente por determinar|Indeterminada|no
134198009|_SUG_Etiologia|perfil probablemente a estudio|Indeterminada|no
134198009|_SUG_Etiologia|perfil probablemente no determinada|Indeterminada|no
134198009|_SUG_Etiologia|perfil probablemente por determinar|Indeterminada|no
134198009|_SUG_Etiologia|por determinar|Indeterminada|no
134198009|_SUG_Etiologia|causa indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|causa indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|causa posiblemente indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|causa posiblemente indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|causa probablemente indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|causa probablemente indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|de origen indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|de origen indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|de origen posiblemente indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|de origen posiblemente indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|de origen probablemente indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|de origen probablemente indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|etiologia indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|etiologia indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|etiologia posiblemente indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|etiologia posiblemente indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|etiologia probablemente indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|etiologia probablemente indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|origen indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|origen indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|origen posiblemente indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|origen posiblemente indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|origen probablemente indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|origen probablemente indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|perfil indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|perfil indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|perfil posiblemente indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|perfil posiblemente indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|perfil probablemente indeterminado de causa doble|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|perfil probablemente indeterminado por doble causa|Indeterminado de causa doble|no
134198009|_SUG_Etiologia|causa con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa posiblemente con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa posiblemente indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa posiblemente indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa posiblemente indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa posiblemente indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa posiblemente pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa posiblemente pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa probablemente con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa probablemente indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa probablemente indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa probablemente indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa probablemente indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa probablemente pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa probablemente pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen posiblemente con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen posiblemente indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen posiblemente indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen posiblemente indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen posiblemente indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen posiblemente pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen posiblemente pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen probablemente con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen probablemente indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen probablemente indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen probablemente indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen probablemente indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen probablemente pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|de origen probablemente pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia posiblemente con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia posiblemente indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia posiblemente indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia posiblemente indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia posiblemente indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia posiblemente pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia posiblemente pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia probablemente con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia probablemente indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia probablemente indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia probablemente indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia probablemente indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia probablemente pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|etiologia probablemente pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen posiblemente con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen posiblemente indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen posiblemente indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen posiblemente indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen posiblemente indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen posiblemente pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen posiblemente pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen probablemente con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen probablemente indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen probablemente indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen probablemente indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen probablemente indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen probablemente pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|origen probablemente pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil posiblemente con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil posiblemente indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil posiblemente indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil posiblemente indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil posiblemente indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil posiblemente pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil posiblemente pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil probablemente con estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil probablemente indeterminada per estudi incomplet|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil probablemente indeterminado (estudio incompleto)|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil probablemente indeterminado pendiente de estudio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil probablemente indeterminado por estudio incompleto|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil probablemente pendent de completar l'estudi|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|perfil probablemente pendent de filiacio|Indeterminado por estudio incompleto|no
134198009|_SUG_Etiologia|causa criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|causa esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|causa indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|causa posiblemente criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|causa posiblemente esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|causa posiblemente indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|causa probablemente criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|causa probablemente esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|causa probablemente indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|de origen criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|de origen esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|de origen indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|de origen posiblemente criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|de origen posiblemente esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|de origen posiblemente indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|de origen probablemente criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|de origen probablemente esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|de origen probablemente indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|etiologia criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|etiologia esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|etiologia indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|etiologia posiblemente criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|etiologia posiblemente esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|etiologia posiblemente indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|etiologia probablemente criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|etiologia probablemente esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|etiologia probablemente indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|origen criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|origen esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|origen indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|origen posiblemente criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|origen posiblemente esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|origen posiblemente indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|origen probablemente criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|origen probablemente esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|origen probablemente indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|perfil criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|perfil esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|perfil indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|perfil posiblemente criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|perfil posiblemente esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|perfil posiblemente indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|perfil probablemente criptogenico|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|perfil probablemente esus|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|perfil probablemente indeterminado|Indeterminado/ESUS|no
134198009|_SUG_Etiologia|causa infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|causa inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|causa insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|causa posiblemente infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|causa posiblemente inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|causa posiblemente insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|causa probablemente infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|causa probablemente inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|causa probablemente insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|de origen infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|de origen inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|de origen insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|de origen posiblemente infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|de origen posiblemente inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|de origen posiblemente insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|de origen probablemente infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|de origen probablemente inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|de origen probablemente insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|etiologia infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|etiologia inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|etiologia insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|etiologia posiblemente infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|etiologia posiblemente inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|etiologia posiblemente insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|etiologia probablemente infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|etiologia probablemente inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|etiologia probablemente insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|origen infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|origen inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|origen insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|origen posiblemente infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|origen posiblemente inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|origen posiblemente insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|origen probablemente infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|origen probablemente inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|origen probablemente insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|perfil infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|perfil inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|perfil insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|perfil posiblemente infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|perfil posiblemente inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|perfil posiblemente insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|perfil probablemente infrecuente|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|perfil probablemente inhabitual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|perfil probablemente insual|Inhabitual o infrecuente|no
134198009|_SUG_Etiologia|causa lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|causa microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|causa posiblemente lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|causa posiblemente microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|causa probablemente lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|causa probablemente microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|de origen lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|de origen microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|de origen posiblemente lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|de origen posiblemente microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|de origen probablemente lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|de origen probablemente microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|etiologia lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|etiologia microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|etiologia posiblemente lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|etiologia posiblemente microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|etiologia probablemente lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|etiologia probablemente microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|origen lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|origen microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|origen posiblemente lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|origen posiblemente microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|origen probablemente lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|origen probablemente microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|perfil lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|perfil microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|perfil posiblemente lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|perfil posiblemente microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|perfil probablemente lacunar|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|perfil probablemente microangiopatica|Lacunar (o microangiopática)|no
134198009|_SUG_Etiologia|causa cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa posiblemente cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa posiblemente diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa posiblemente malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa posiblemente secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa posiblemente secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa probablemente cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa probablemente diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa probablemente malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa probablemente secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa probablemente secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen posiblemente cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen posiblemente diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen posiblemente malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen posiblemente secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen posiblemente secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen probablemente cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen probablemente diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen probablemente malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen probablemente secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen probablemente secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|de origen secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia posiblemente cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia posiblemente diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia posiblemente malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia posiblemente secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia posiblemente secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia probablemente cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia probablemente diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia probablemente malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia probablemente secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia probablemente secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|etiologia secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen posiblemente cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen posiblemente diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen posiblemente malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen posiblemente secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen posiblemente secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen probablemente cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen probablemente diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen probablemente malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen probablemente secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen probablemente secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|origen secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil posiblemente cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil posiblemente diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil posiblemente malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil posiblemente secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil posiblemente secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil probablemente cavernoma de circunvolucion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil probablemente diseccio|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil probablemente malformacion arteriovenosa|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil probablemente secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil probablemente secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|perfil secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|secundaria a diseccion|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|secundaria a malformacion vascular|Secundaria a malformación vascular/aneurisma|no
134198009|_SUG_Etiologia|causa posiblemente secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|causa probablemente secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|causa secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|de origen posiblemente secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|de origen probablemente secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|de origen secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|etiologia posiblemente secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|etiologia probablemente secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|etiologia secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|origen posiblemente secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|origen probablemente secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|origen secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|perfil posiblemente secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|perfil probablemente secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|perfil secundaria a tumor|Secundaria a tumor|no
134198009|_SUG_Etiologia|secundaria a tumor|Secundaria a tumor|no
1386000|_SUG_Hemorragia_cerebral|acv hemorragia|Hemorragia cerebral|no
1386000|_SUG_Hemorragia_cerebral|avc hemorragia|Hemorragia cerebral|no
1386000|_SUG_Hemorragia_cerebral|hematoma|Hemorragia cerebral|no
1386000|_SUG_Hemorragia_cerebral|hematoma cerebral|Hemorragia cerebral|no
1386000|_SUG_Hemorragia_cerebral|hematoma intracraneal|Hemorragia cerebral|no
1386000|_SUG_Hemorragia_cerebral|hematoma intraparenquimatoso|Hemorragia cerebral|no
1386000|_SUG_Hemorragia_cerebral|hematoma parenquimatoso|Hemorragia cerebral|no
1386000|_SUG_Hemorragia_cerebral|hemorragia|Hemorragia cerebral|no
1386000|_SUG_Hemorragia_cerebral|hemorragia cerebral|Hemorragia cerebral|no
1386000|_SUG_Hemorragia_cerebral|hemorragia intracerebral|Hemorragia cerebral|no
1386000|_SUG_Hemorragia_cerebral|hemorragia parenquimatosa|Hemorragia cerebral|no
1386000|_SUG_Hemorragia_cerebral|hemorragia parenquimatosa cerebral masiva|Hemorragia cerebral|no
1386000|_SUG_Hemorragia_cerebral|hic|Hemorragia cerebral|no
1386000|_SUG_Hemorragia_cerebral|ictus hemorragia|Hemorragia cerebral|no
422504002|_SUG_Ictus_isquemico|avc isquemia|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|e. cerebrovascular aguda isquemia: infarto|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|ecva isquemia|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|ecva isquemia: infarto|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|ecva isquemia: infarto cerebral|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|ecva: infartos isquemicos|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|enfermedad cerebrovascular aguda isquemia|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|ictus|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|ictus isquemia|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|ictus isquemia agudo|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|ictus isquemia con transformacion hemorragia|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|infarto|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|infarto agudo|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|infarto cerebeloso|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|infarto cerebral|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|infarto isquemia|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|infarto isquemia agudo|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|infarto isquemia cerebral|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|infarto isquemicos|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|isquemia en territorio cortical|Ictus isquémico|no
422504002|_SUG_Ictus_isquemico|transformacion hemorragia|Otros|no
422504002|_SUG_Ictus_isquemico|sufusion hemorragia|Otros|no
422504002|_SUG_Ictus_isquemico|accidente cerebrovascular|Otros|no
422504002|_SUG_Ictus_isquemico|avc|Otros|no
422504002|_SUG_Ictus_isquemico|sindrome de alarma capsular|Otros|no
422504002|_SUG_Ictus_isquemico|sindrome sensitivo motor|Otros|no
422504002|_SUG_Ictus_isquemico|sindrome sensitivo-motor regresivo|Otros|no
00000019|_SUG_Lateralizacion|ambas|Bilateral|no
00000019|_SUG_Lateralizacion|bihemisferico|Bilateral|no
00000019|_SUG_Lateralizacion|bilaterales|Bilateral|no
00000019|_SUG_Lateralizacion|D|Derecha|no
00000019|_SUG_Lateralizacion|dcha|Derecha|no
00000019|_SUG_Lateralizacion|dcho|Derecha|no
00000019|_SUG_Lateralizacion|derecho|Derecha|no
00000019|_SUG_Lateralizacion|dret|Derecha|no
00000019|_SUG_Lateralizacion|dreta|Derecha|no
00000019|_SUG_Lateralizacion|E|Izquierda|no
00000019|_SUG_Lateralizacion|e|Izquierda|no
00000019|_SUG_Lateralizacion|esq|Izquierda|no
00000019|_SUG_Lateralizacion|esq.|Izquierda|no
00000019|_SUG_Lateralizacion|esquerre|Izquierda|no
00000019|_SUG_Lateralizacion|I|Izquierda|no
00000019|_SUG_Lateralizacion|izda|Izquierda|no
00000019|_SUG_Lateralizacion|izdo|Izquierda|no
00000019|_SUG_Lateralizacion|izq|Izquierda|no
00000019|_SUG_Lateralizacion|izquierda|Izquierda|no
00000019|_SUG_Lateralizacion|tronco cerebral|Tronco cerebral|no
246267002|_SUG_Localizacion|bulbar|Bulbar|no
246267002|_SUG_Localizacion|cerebelosa|Cerebelosa|no
246267002|_SUG_Localizacion|cortical|Cortical|no
246267002|_SUG_Localizacion|fronto insular|Frontal|no
246267002|_SUG_Localizacion|fronto|Frontal y occipital|no
246267002|_SUG_Localizacion|fronto occipital|Frontal y occipital|no
246267002|_SUG_Localizacion|fronto y occipital|Frontal y occipital|no
246267002|_SUG_Localizacion|fronto temporo insular|Frontal y temporal|no
246267002|_SUG_Localizacion|indeterminado|Indeterminada|no
246267002|_SUG_Localizacion|parcial|Indeterminada|no
246267002|_SUG_Localizacion|territorio indeterminado|Indeterminada|no
246267002|_SUG_Localizacion|poci|Infarto de circulación posterior o POCI|no
246267002|_SUG_Localizacion|infarto lacunar|Infarto lacunar o LACI|no
246267002|_SUG_Localizacion|laci|Infarto lacunar o LACI|no
246267002|_SUG_Localizacion|lacunar|Infarto lacunar o LACI|no
246267002|_SUG_Localizacion|infarto parcial de circulacion anterior|Infarto parcial de circulación anterior o PACI|no
246267002|_SUG_Localizacion|paci|Infarto parcial de circulación anterior o PACI|no
246267002|_SUG_Localizacion|infarto total de circulacion anterior|Infarto total de circulación anterior o TACI|no
246267002|_SUG_Localizacion|taci|Infarto total de circulación anterior o TACI|no
246267002|_SUG_Localizacion|intraventricular|Intraventricular|no
246267002|_SUG_Localizacion|ventriculos|Intraventricular|no
246267002|_SUG_Localizacion|lobar|Lobar|no
246267002|_SUG_Localizacion|occipital|Occipital|no
246267002|_SUG_Localizacion|parietal|Parietal|no
246267002|_SUG_Localizacion|parietooccipital|Parietal y occipital|no
246267002|_SUG_Localizacion|infarto de circulacion posterior|Posterior|no
246267002|_SUG_Localizacion|posterior|Posterior|no
246267002|_SUG_Localizacion|protuberancial|Posterior|no
246267002|_SUG_Localizacion|basilar|Posterior/tronco/bulbar|no
246267002|_SUG_Localizacion|capsulo talamic|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|caudado|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|corona radiada|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|ganglicapsular|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|ganglios basales|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|ganglios de la base|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|ggbb|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|lenticular|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|lenticular capsular|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|lenticular capsulotalamico|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|palido|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|profunda|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|profundes|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|putamen|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|putaminal|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|talamica|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|talamo|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|talamo capuslar|Profunda o ganglios de la base|no
246267002|_SUG_Localizacion|subcorticals|Subcortical|no
246267002|_SUG_Localizacion|emporo insular|Temporal|no
246267002|_SUG_Localizacion|temporal|Temporal|no
246267002|_SUG_Localizacion|temporal basal|Temporal y profunda|no
246267002|_SUG_Localizacion|tronco|Troncal|no
273729003|_SUG_mRankin|escala de rankin modificada 0|mRankin|no
273729003|_SUG_mRankin|mrankin 0|mRankin|no
273729003|_SUG_mRankin|mrankinscale 0|mRankin|no
273729003|_SUG_mRankin|mrs 0|mRankin|no
273729003|_SUG_mRankin|rankin 0|mRankin|no
450741005|_SUG_NIHSS|0 en la escala nihss|NIHSS|no
450741005|_SUG_NIHSS|escala nihss 0|NIHSS|no
450741005|_SUG_NIHSS|escala nihss es de 0 puntos|NIHSS|no
450741005|_SUG_NIHSS|nhiss 0|NIHSS|no
450741005|_SUG_NIHSS|nih 0|NIHSS|no
450741005|_SUG_NIHSS|nihaa 0|NIHSS|no
450741005|_SUG_NIHSS|nihss 0|NIHSS|no
450741005|_SUG_NIHSS|nishss 0|NIHSS|no
450741005|_SUG_NIHSS|nissh 0|NIHSS|no
450741005|_SUG_NIHSS|puntuacion total nih:0|NIHSS|no
00000025|_SUG_Puerta_aguja|puerta aguja|Tiempo puerta-aguja|no
00000024|_SUG_Recanalizacion|recanalizacion|Recanalización|no
34227000|_SUG_TAC_craneal|tc arterias cerebrales|Angiotomografía computarizada|no
34227000|_SUG_TAC_craneal|tac|TAC|no
34227000|_SUG_TAC_craneal|tc|TAC|no
34227000|_SUG_TAC_craneal|tac - craneal|Tac craneal|no
34227000|_SUG_TAC_craneal|tac cerebral|Tac craneal|no
34227000|_SUG_TAC_craneal|tac cerebro|Tac craneal|no
34227000|_SUG_TAC_craneal|tac craneal|Tac craneal|no
34227000|_SUG_TAC_craneal|tac craneo|Tac craneal|no
34227000|_SUG_TAC_craneal|tac crani|Tac craneal|no
34227000|_SUG_TAC_craneal|tac crani al|Tac craneal|no
34227000|_SUG_TAC_craneal|tac cranial|Tac craneal|no
34227000|_SUG_TAC_craneal|tac de cap|Tac craneal|no
34227000|_SUG_TAC_craneal|tac de craneo|Tac craneal|no
34227000|_SUG_TAC_craneal|tacs craneales|Tac craneal|no
34227000|_SUG_TAC_craneal|tc - craneal|Tac craneal|no
34227000|_SUG_TAC_craneal|tc cerebral|Tac craneal|no
34227000|_SUG_TAC_craneal|tc cerebro|Tac craneal|no
34227000|_SUG_TAC_craneal|tc craneal|Tac craneal|no
34227000|_SUG_TAC_craneal|tc crani|Tac craneal|no
34227000|_SUG_TAC_craneal|tc crani al|Tac craneal|no
34227000|_SUG_TAC_craneal|tc cranial|Tac craneal|no
34227000|_SUG_TAC_craneal|tc de cap|Tac craneal|no
34227000|_SUG_TAC_craneal|tc de craneo|Tac craneal|no
34227000|_SUG_TAC_craneal|tomografia axial computeritzada de cap|Tac craneal|no
34227000|_SUG_TAC_craneal|tomografia de cap|Tac craneal|no
34227000|_SUG_TAC_craneal|tac perfusion cerebral|TAC-perfusión|no
34227000|_SUG_TAC_craneal|tac perfusioncerebral|TAC-perfusión|no
34227000|_SUG_TAC_craneal|tc perfusion cerebral|TAC-perfusión|no
34227000|_SUG_TAC_craneal|tc perfusioncerebral|TAC-perfusión|no
00000008|_SUG_Test_de_disfagia|prueba de disfagia|Test de disfagia|no
00000007|_SUG_Test_de_disfagia|test de deglucion|Test de disfagia|no
00000007|_SUG_Test_de_disfagia|test de disfagia|Test de disfagia|no
00000007|_SUG_Test_de_disfagia|test deglucion|Test de disfagia|no
00000007|_SUG_Test_de_disfagia|test mecv-v|Test de disfagia|no
108972005|_SUG_Tratamiento_antiagregante|a.a.s.|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|aas|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|abciximab|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|ac acetilsalicilico|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|acetil salicilic-acid|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|acetilsalicilico|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|acetilsalicilico acido|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|acetylsalicylic acid|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|acido acetilsalicilico|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|adiro|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|agrastat|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|aspirina|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|brilique|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|cangrelor|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|cilostazol|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|clopidogrel|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|combinations|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|dipyridamole|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|disgren|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|duoplavin|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|ekistol|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|hepraina|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|persantin|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|plavix|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|pletal|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|prasugler|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|reopro|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|ticagrelor|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|ticlopidine|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|tiklid|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|tirofiban|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|triflusal|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|tromalyt|Tratamiento antiagregante|no
108972005|_SUG_Tratamiento_antiagregante|vatoud|Tratamiento antiagregante|no
81839001|_SUG_Tratamiento_anticoagulante|acenocumarol|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|aldocumar|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|apixaban|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|bemiparin|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|clexane|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|dabigatran|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|dabigatran etexilate|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|dalteparin|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|edoxaban|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|eliquis|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|enoxaparin|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|fragmin|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|fraxiparina|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|hbpm|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|heparin|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|heparina|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|hibor|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|innohep|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|lixiana|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|nadroparin|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|parnaparin|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|pradaxa|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|reviparin|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|rivaroxaban|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|sintrom|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|warfarin|Tratamiento anticoagulante|no
81839001|_SUG_Tratamiento_anticoagulante|xarelto|Tratamiento anticoagulante|no
433112001|_SUG_Trombectomia_mecanica|angioradiologia intervencionista|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|arteriografia trombectomia|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|embolectomia mecanica|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|procedimiento de revascularizacion|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|reperfusion intraateria|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|rescate endovascular|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|rescate intraarterial|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|terapia de reperfusion|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|terapia de rescate|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|terapia endovascular|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|terapia endovascular (trombectomia mecanica)|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tev|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tev (trombectomia mecanica)|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tev mecanica|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tractament intraarterial|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tractament mecanic endovascular|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tractament neurovascular|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento agudo mecanico|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento de reperfusion|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento de reperfusion intrarterial|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento de reperfusionmediante trombectomia mecanica|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento de repermeabilizacion|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento de rescate|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento de revascularizacion|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento de revascularizacion intraarterial|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento endovascular|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento endovascular mediante trombectomia mecnica|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento intraarterial|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento intraarterial primario|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento mecanico del ictus|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento neurointervencionista|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento recanalizador|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento recanalizador endovenoso|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento reperfusion|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento rescate endovascular|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tratamiento revascularizador|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomia|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomia cerebrala|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomia endovascular|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomia endovenosa|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomia extra e intracraneal mecanica|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomia intra i extra craneal mecanica|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomia intra y extracranea|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomia intracraneal|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomia intracraneal mecanica|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomia mecanica|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomia mecanica endovascular|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomia mecanica primaria|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomia trombectomiamecanica|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomiacerebrala|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|trombectomiamecanica|trombectomía mecánica|no
433112001|_SUG_Trombectomia_mecanica|tto endovascular|trombectomía mecánica|no
00000006|_SUG_Trombolisis_intraarterial|trombolisis ia|trombólisis intraarterial|no
00000006|_SUG_Trombolisis_intraarterial|trombolisis intraarterial|trombólisis intraarterial|no
472191000119101|_SUG_Trombolisis_intravenosa|actylise|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|ecas iv|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolisi amb rtpa ev|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolisis|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolisis con alteplase|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolisis con r-tpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolisis con rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolisis con rtpa endovenoso|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolisis con rtpa intravenosa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolisis endovenosa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolisis endovenosa con rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolisis endovenosa rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolisis ev con rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolisis iv|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolisis rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolisis sistemica con rtpa ev|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolitico|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolitico amb rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolitico con rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|fibrinolizado|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|procedimiento de revascularizacion|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|rtpa ev|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|rtpaev|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tecneplasa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|terapia de reperfusion|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|terapia de rescate|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tnk|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tpa ev|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tractament amb rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tractament amb rtpa endovenos|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tractament endovenos|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tractament fibrinolitic ev|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tractament fibrinolitic|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tractament fibrinolitic|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tractament fibrinolitic endovenos amb rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tractament rpta ev|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tractat amb firbinolisi|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento con alteplasa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento con fibrinolisis ev|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento con rt-pa intravenoso|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento con rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento con rtpa ev|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento de repefusion cerebral con r-tpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento de reperfusion|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento de reperfusion aguda mendiante fibrinolisis ev|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento de reperfusion con fibrinolisis|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento de reperfusion con fibrinolisis ev|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento de reperfusion con rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento de reperfusion de rpta endovenoso|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento de reperfusion en fase aguda con rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento de reperfusion ev|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento de repermeabilizacion|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento de revascularizacion|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento endovenoso|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento fibrinolitico|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento fibrinolitico con alteplase|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento fibrinolitico con rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento fibrinolitico con rtpa endovenosa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento fibrinolitico con rtpa ev|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento fibrinolitico endovenoso|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento fibrinolitico ev con rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento fibrinolitico rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento fibrinolotico iv|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento recanalizador|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento recanalizador con fibrinolisis iv|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento recanalizador endovenoso|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento reperfusion|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento reperfusor con fibrinolitico endovenoso|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento reperfusor endovenoso|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento revascularizador|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento trombolitico|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento trombolitico con rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento trombolitico con tpa endovenoso|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento trombolitico intravenoso|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento trombolitico intravenoso con rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tratamiento trombolitico rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|trombolisado|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|trombolisis|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|trombolisis cerebral|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|trombolisis endovenosa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|trombolisis ev|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|trombolisis intravenosa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|trombolisis sistemica endovenosa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|trombolisisendovenosa con rtpa|Trombólisis intravenosa|no
472191000119101|_SUG_Trombolisis_intravenosa|tto trombolitico con rtpa|Trombólisis intravenosa|no
