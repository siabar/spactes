C0000001|_SUG_Ictus_isquemico|accidente cerebrovascular
C0000001|_SUG_Ictus_isquemico|AVC
C0000001|_SUG_Ictus_isquemico|AVC isquemic
C0000001|_SUG_Ictus_isquemico|ECVA ISQUEMICA
C0000001|_SUG_Ictus_isquemico|ECVA ISQUEMICA: INFARTO
C0000001|_SUG_Ictus_isquemico|ECVA: INFARTOS ISQUEMICOS
C0000001|_SUG_Ictus_isquemico|ictus
C0000001|_SUG_Ictus_isquemico|ICTUS ISQUEMIC
C0000001|_SUG_Ictus_isquemico|ictus isquemico con transformacion hemorragica
C0000001|_SUG_Ictus_isquemico|Infart isquemic
C0000001|_SUG_Ictus_isquemico|Infart
C0000001|_SUG_Ictus_isquemico|Infartos
C0000001|_SUG_Ictus_isquemico|Infartos isquemicos
C0000001|_SUG_Ictus_isquemico|infarto
C0000001|_SUG_Ictus_isquemico|infarto cerebral
C0000001|_SUG_Ictus_isquemico|infarto isquemico
C0000001|_SUG_Ictus_isquemico|Infarto isquemico agudo
C0000001|_SUG_Ictus_isquemico|sufusion hemorragica
C0000001|_SUG_Ictus_isquemico|transformacion hemorragica
C0000002|_SUG_Ataque_isquemico_transitorio|ACCIDENTE TRANSITORI ISQUEMICO
C0000002|_SUG_Ataque_isquemico_transitorio|AIT
C0000002|_SUG_Ataque_isquemico_transitorio|ataque isquemico transitorio
C0000002|_SUG_Ataque_isquemico_transitorio|ICTUS MINOR
C0000002|_SUG_Ataque_isquemico_transitorio|Infarto clinicamente regresivo
C0000002|_SUG_Ataque_isquemico_transitorio|Sindrome sensitivo-motor regresivo
C0000002|_SUG_Ataque_isquemico_transitorio|TIA
C0000003|_SUG_Hemorragia_cerebral|AVC HEMORRAGIC
C0000003|_SUG_Hemorragia_cerebral|HEMATOMA
C0000003|_SUG_Hemorragia_cerebral|hematoma cerebral
C0000003|_SUG_Hemorragia_cerebral|HEMORRAGIA
C0000003|_SUG_Hemorragia_cerebral|hemorragia cerebral
C0000003|_SUG_Hemorragia_cerebral|hemorragia intracerebral
C0000003|_SUG_Hemorragia_cerebral|HEMORRAGIA PARENQUIMATOSA CEREBRAL MASIVA
C0000003|_SUG_Hemorragia_cerebral|ictus hemorragico
C0000004|_SUG_Trombolisis_intravenosa|ECAS IV
C0000004|_SUG_Trombolisis_intravenosa|fibrinolotico
C0000004|_SUG_Trombolisis_intravenosa|fibrinolisis
C0000004|_SUG_Trombolisis_intravenosa|fibrinolisis endovenosa
C0000004|_SUG_Trombolisis_intravenosa|fibrinolisis iv
C0000004|_SUG_Trombolisis_intravenosa|fibrinolisis sistemica con rtPA ev
C0000004|_SUG_Trombolisis_intravenosa|rtPA
C0000004|_SUG_Trombolisis_intravenosa|tPAev
C0000004|_SUG_Trombolisis_intravenosa|tractat amb firbinolisi
C0000004|_SUG_Trombolisis_intravenosa|trombolisis
C0000004|_SUG_Trombolisis_intravenosa|tratamiento con alteplasa
C0000004|_SUG_Trombolisis_intravenosa|Tratamiento con RTPA
C0000004|_SUG_Trombolisis_intravenosa|tratamiento fibrinolitico
C0000004|_SUG_Trombolisis_intravenosa|tratamiento trombolitico
C0000004|_SUG_Trombolisis_intravenosa|trombolisis intravenosa
C0000005|_SUG_Trombectomia_mecanica|TEV
C0000005|_SUG_Trombectomia_mecanica|trombectomia
C0000005|_SUG_Trombectomia_mecanica|tratamiento agudo mecanico
C0000005|_SUG_Trombectomia_mecanica|tratamiento endovascular
C0000005|_SUG_Trombectomia_mecanica|Trombectomia endovascular
C0000005|_SUG_Trombectomia_mecanica|Trombectomia mecanica
C0000006|_SUG_Trombolisis_intraarterial|trombolisis ia
C0000006|_SUG_Trombolisis_intraarterial|trombolisis intraarterial
C0000007|_SUG_Test_de_disfagia|test de deglucion
C0000007|_SUG_Test_de_disfagia|test de disfagia
C0000011|_SUG_mRankin|Escala de Rankin modificada 0
C0000012|_SUG_NIHSS|escala NIHSS es de 0 puntos
C0000012|_SUG_NIHSS|Escala NIHSS 0
C0000012|_SUG_NIHSS|PUNTUACION TOTAL NIH:0
C0000010|_SUG_ASPECTS|ASPECTS 0
C0000010|_SUG_ASPECTS|ASPECTS score 0
C0000011|_SUG_mRankin|mRankinScale 0
C0000011|_SUG_mRankin|mRankin 0
C0000011|_SUG_mRankin|mRS 0
C0000011|_SUG_mRankin|Rankin 0
C0000012|_SUG_NIHSS|NIH 0
C0000012|_SUG_NIHSS|NIHSS 0
C0000012|_SUG_NIHSS|NHISS 0
C0000012|_SUG_NIHSS|NISHSS 0
C0000012|_SUG_NIHSS|NISSH 0
C0000013|_SUG_Tratamiento_anticoagulante|acenocumarol
C0000013|_SUG_Tratamiento_anticoagulante|aldocumar
C0000013|_SUG_Tratamiento_anticoagulante|apixaban
C0000013|_SUG_Tratamiento_anticoagulante|B01AA03
C0000013|_SUG_Tratamiento_anticoagulante|B01AA07
C0000013|_SUG_Tratamiento_anticoagulante|B01AB01
C0000013|_SUG_Tratamiento_anticoagulante|B01AB04
C0000013|_SUG_Tratamiento_anticoagulante|B01AB05
C0000013|_SUG_Tratamiento_anticoagulante|B01AB06
C0000013|_SUG_Tratamiento_anticoagulante|B01AB07
C0000013|_SUG_Tratamiento_anticoagulante|B01AB08
C0000013|_SUG_Tratamiento_anticoagulante|B01AB12
C0000013|_SUG_Tratamiento_anticoagulante|B01AE07
C0000013|_SUG_Tratamiento_anticoagulante|B01AF01
C0000013|_SUG_Tratamiento_anticoagulante|B01AF02
C0000013|_SUG_Tratamiento_anticoagulante|B01AF03
C0000013|_SUG_Tratamiento_anticoagulante|bemiparin
C0000013|_SUG_Tratamiento_anticoagulante|clexane
C0000013|_SUG_Tratamiento_anticoagulante|Dabigatran
C0000013|_SUG_Tratamiento_anticoagulante|dabigatran etexilate
C0000013|_SUG_Tratamiento_anticoagulante|dalteparin
C0000013|_SUG_Tratamiento_anticoagulante|edoxaban
C0000013|_SUG_Tratamiento_anticoagulante|eliquis
C0000013|_SUG_Tratamiento_anticoagulante|enoxaparin
C0000013|_SUG_Tratamiento_anticoagulante|fragmin
C0000013|_SUG_Tratamiento_anticoagulante|fraxiparina
C0000013|_SUG_Tratamiento_anticoagulante|heparin
C0000013|_SUG_Tratamiento_anticoagulante|Heparina
C0000013|_SUG_Tratamiento_anticoagulante|hibor
C0000013|_SUG_Tratamiento_anticoagulante|lixiana
C0000013|_SUG_Tratamiento_anticoagulante|nadroparin
C0000013|_SUG_Tratamiento_anticoagulante|parnaparin
C0000013|_SUG_Tratamiento_anticoagulante|pradaxa
C0000013|_SUG_Tratamiento_anticoagulante|reviparin
C0000013|_SUG_Tratamiento_anticoagulante|rivaroxaban
C0000013|_SUG_Tratamiento_anticoagulante|sintrom
C0000013|_SUG_Tratamiento_anticoagulante|warfarin
C0000013|_SUG_Tratamiento_anticoagulante|xarelto
C0000016|_SUG_Tratamiento_antiagregante|AAS
C0000016|_SUG_Tratamiento_antiagregante|abciximab
C0000016|_SUG_Tratamiento_antiagregante|AC ACETILSALICILICO
C0000016|_SUG_Tratamiento_antiagregante|acetylsalicylic acid
C0000016|_SUG_Tratamiento_antiagregante|acetylsalicylic acid, combinations with proton pump inhibitors
C0000016|_SUG_Tratamiento_antiagregante|Acido acetilsalicilico
C0000016|_SUG_Tratamiento_antiagregante|Adiro
C0000016|_SUG_Tratamiento_antiagregante|agrastat
C0000016|_SUG_Tratamiento_antiagregante|Aspirina
C0000016|_SUG_Tratamiento_antiagregante|B01AC04
C0000016|_SUG_Tratamiento_antiagregante|B01AC05
C0000016|_SUG_Tratamiento_antiagregante|B01AC06
C0000016|_SUG_Tratamiento_antiagregante|B01AC07
C0000016|_SUG_Tratamiento_antiagregante|B01AC13
C0000016|_SUG_Tratamiento_antiagregante|B01AC17
C0000016|_SUG_Tratamiento_antiagregante|B01AC18
C0000016|_SUG_Tratamiento_antiagregante|B01AC22
C0000016|_SUG_Tratamiento_antiagregante|B01AC23
C0000016|_SUG_Tratamiento_antiagregante|B01AC24
C0000016|_SUG_Tratamiento_antiagregante|B01AC25
C0000016|_SUG_Tratamiento_antiagregante|B01AC30
C0000016|_SUG_Tratamiento_antiagregante|B01AC56
C0000016|_SUG_Tratamiento_antiagregante|brilique
C0000016|_SUG_Tratamiento_antiagregante|cangrelor
C0000016|_SUG_Tratamiento_antiagregante|cido acetilsalicilico
C0000016|_SUG_Tratamiento_antiagregante|cilostazol
C0000016|_SUG_Tratamiento_antiagregante|clopidogrel
C0000016|_SUG_Tratamiento_antiagregante|combinations
C0000016|_SUG_Tratamiento_antiagregante|dipyridamole
C0000016|_SUG_Tratamiento_antiagregante|disgren
C0000016|_SUG_Tratamiento_antiagregante|ekistol
C0000016|_SUG_Tratamiento_antiagregante|persantin
C0000016|_SUG_Tratamiento_antiagregante|plavix
C0000016|_SUG_Tratamiento_antiagregante|pletal
C0000016|_SUG_Tratamiento_antiagregante|prasugler
C0000016|_SUG_Tratamiento_antiagregante|reopro
C0000016|_SUG_Tratamiento_antiagregante|ticagrelor
C0000016|_SUG_Tratamiento_antiagregante|ticlopidine
C0000016|_SUG_Tratamiento_antiagregante|tiklid
C0000016|_SUG_Tratamiento_antiagregante|tirofiban
C0000016|_SUG_Tratamiento_antiagregante|triflusal
C0000017|_SUG_Arteria_afectada|A.COROIDEA ANT
C0000017|_SUG_Arteria_afectada|A2
C0000017|_SUG_Arteria_afectada|AB
C0000017|_SUG_Arteria_afectada|ACA
C0000017|_SUG_Arteria_afectada|ACC
C0000017|_SUG_Arteria_afectada|ACI
C0000017|_SUG_Arteria_afectada|ACI-T
C0000017|_SUG_Arteria_afectada|ACM
C0000017|_SUG_Arteria_afectada|ACP
C0000017|_SUG_Arteria_afectada|ACS
C0000017|_SUG_Arteria_afectada|AICA
C0000017|_SUG_Arteria_afectada|art Vertebral
C0000017|_SUG_Arteria_afectada|Arteria basilar
C0000017|_SUG_Arteria_afectada|Arteria carotida comun
C0000017|_SUG_Arteria_afectada|Arteria carotida interna
C0000017|_SUG_Arteria_afectada|Arteria carotida interna terminal
C0000017|_SUG_Arteria_afectada|arteria carotide
C0000017|_SUG_Arteria_afectada|Arteria cerebelosa anteroinferior
C0000017|_SUG_Arteria_afectada|Arteria cerebelosa posteroinferior
C0000017|_SUG_Arteria_afectada|Arteria cerebelosa superior
C0000017|_SUG_Arteria_afectada|Arteria cerebral anterior
C0000017|_SUG_Arteria_afectada|Arteria cerebral media
C0000017|_SUG_Arteria_afectada|Arteria cerebral media segmento
C0000017|_SUG_Arteria_afectada|arteria cerebral mitja
C0000017|_SUG_Arteria_afectada|Arteria cerebral posterior
C0000017|_SUG_Arteria_afectada|Arteria coroidea anterior
C0000017|_SUG_Arteria_afectada|Arteria coroidea posterior
C0000017|_SUG_Arteria_afectada|Arteria lenticuloestriada
C0000017|_SUG_Arteria_afectada|Arteria vertebral
C0000017|_SUG_Arteria_afectada|ARTERIES CEREBRALS MITGES
C0000017|_SUG_Arteria_afectada|C1
C0000017|_SUG_Arteria_afectada|carotida primitiva
C0000017|_SUG_Arteria_afectada|carotidea
C0000017|_SUG_Arteria_afectada|CAROTIDEA
C0000017|_SUG_Arteria_afectada|INDETERM I NA DO
C0000017|_SUG_Arteria_afectada|indeterminado
C0000017|_SUG_Arteria_afectada|M1
C0000017|_SUG_Arteria_afectada|M6
C0000017|_SUG_Arteria_afectada|M2
C0000017|_SUG_Arteria_afectada|M3
C0000017|_SUG_Arteria_afectada|M4
C0000017|_SUG_Arteria_afectada|M5
C0000017|_SUG_Arteria_afectada|nucleo lenticular
C0000017|_SUG_Arteria_afectada|PICA
C0000017|_SUG_Arteria_afectada|territorio indeterminado
C0000017|_SUG_Arteria_afectada|TICA
C0000017|_SUG_Arteria_afectada|V1
C0000017|_SUG_Arteria_afectada|VB
C0000017|_SUG_Arteria_afectada|VERTEBR BASILAR
C0000017|_SUG_Arteria_afectada|vertebro-basilar
C0000017|_SUG_Arteria_afectada|vertebrobasilar
C0000018|_SUG_Localizacion|BULBAR
C0000018|_SUG_Localizacion|capsulo-talamic
C0000018|_SUG_Localizacion|capsulotalamico
C0000018|_SUG_Localizacion|caudado
C0000018|_SUG_Localizacion|cerebelosa
C0000018|_SUG_Localizacion|corona radiada
C0000018|_SUG_Localizacion|cortical
C0000018|_SUG_Localizacion|frontal
C0000018|_SUG_Localizacion|fronto-insular
C0000018|_SUG_Localizacion|fronto-temporo-insular
C0000018|_SUG_Localizacion|ganglicapsular
C0000018|_SUG_Localizacion|GANGLIOS BASALES
C0000018|_SUG_Localizacion|ganglios de la base
C0000018|_SUG_Localizacion|ggbb
C0000018|_SUG_Localizacion|Infarto de circulacion posterior
C0000018|_SUG_Localizacion|Infarto lacunar
C0000018|_SUG_Localizacion|Infarto parcial de circulacion anterior
C0000018|_SUG_Localizacion|Infarto total de circulacion anterior
C0000018|_SUG_Localizacion|Intraventricular
C0000018|_SUG_Localizacion|LACI
C0000018|_SUG_Localizacion|LACUNAR
C0000018|_SUG_Localizacion|lenticular
C0000018|_SUG_Localizacion|Lobar
C0000018|_SUG_Localizacion|occipital
C0000018|_SUG_Localizacion|PACI
C0000018|_SUG_Localizacion|palido
C0000018|_SUG_Localizacion|parcial
C0000018|_SUG_Localizacion|parietal
C0000018|_SUG_Localizacion|parietooccipital
C0000018|_SUG_Localizacion|POCI
C0000018|_SUG_Localizacion|posterior
C0000018|_SUG_Localizacion|profunda
C0000018|_SUG_Localizacion|profundes
C0000018|_SUG_Localizacion|putamen
C0000018|_SUG_Localizacion|subcorticals
C0000018|_SUG_Localizacion|TACI
C0000018|_SUG_Localizacion|talamica
C0000018|_SUG_Localizacion|talamo
C0000018|_SUG_Localizacion|talamo-capuslar
C0000018|_SUG_Localizacion|temporal
C0000018|_SUG_Localizacion|tronco
C0000018|_SUG_Localizacion|ventriculos
C0000019|_SUG_Lateralizacion|ambas
C0000019|_SUG_Lateralizacion|bilateral
C0000019|_SUG_Lateralizacion|bilaterales
C0000019|_SUG_Lateralizacion|D
C0000019|_SUG_Lateralizacion|Dcha
C0000019|_SUG_Lateralizacion|Derecha
C0000019|_SUG_Lateralizacion|DERECHOS
C0000019|_SUG_Lateralizacion|dret
C0000019|_SUG_Lateralizacion|dreta
C0000019|_SUG_Lateralizacion|E
C0000019|_SUG_Lateralizacion|e
C0000019|_SUG_Lateralizacion|esq
C0000019|_SUG_Lateralizacion|esquerra
C0000019|_SUG_Lateralizacion|esquerres
C0000019|_SUG_Lateralizacion|I
C0000019|_SUG_Lateralizacion|izda
C0000019|_SUG_Lateralizacion|Izq
C0000019|_SUG_Lateralizacion|izquierda
C0000019|_SUG_Lateralizacion|Tronco cerebral
C0000020|_SUG_Etiologia|a estudio
C0000020|_SUG_Etiologia|aneurisma
C0000020|_SUG_Etiologia|angiopatia amiloide
C0000020|_SUG_Etiologia|ateromatosis
C0000020|_SUG_Etiologia|aterosclerotico
C0000020|_SUG_Etiologia|Aterotrombotico
C0000020|_SUG_Etiologia|Cardioembolico
C0000020|_SUG_Etiologia|Cavernoma de circunvolucion
C0000020|_SUG_Etiologia|criptogenico
C0000020|_SUG_Etiologia|Diseccio
C0000020|_SUG_Etiologia|embolico
C0000020|_SUG_Etiologia|ESUS
C0000020|_SUG_Etiologia|Hipertensiva
C0000020|_SUG_Etiologia|indeterminada
C0000020|_SUG_Etiologia|Indeterminado de causa doble
C0000020|_SUG_Etiologia|Indeterminado por estudio incompleto
C0000020|_SUG_Etiologia|infrecuente
C0000020|_SUG_Etiologia|Inhabitual
C0000020|_SUG_Etiologia|Lacunar
C0000020|_SUG_Etiologia|malformacion arteriovenosa
C0000020|_SUG_Etiologia|mecanisme embolic
C0000020|_SUG_Etiologia|secundaria a malformacion vascular
C0000020|_SUG_Etiologia|secundaria a tumor
C0000021|_SUG_TAC_craneal|AgioTAC
C0000021|_SUG_TAC_craneal|TAC
C0000021|_SUG_TAC_craneal|TAC crani al
C0000021|_SUG_TAC_craneal|TAC cerebral
C0000021|_SUG_TAC_craneal|TAC craneal
C0000021|_SUG_TAC_craneal|Tac de craneo
C0000021|_SUG_TAC_craneal|TC
C0000021|_SUG_TAC_craneal|TC craneal
C0000021|_SUG_TAC_craneal|TC cranial
C0000021|_SUG_TAC_craneal|TC de craneo
C0000017|_SUG_Arteria_afectada|A. carotida interna
C0000017|_SUG_Arteria_afectada|ACM-ACA
C0000017|_SUG_Arteria_afectada|Art Basilar
C0000017|_SUG_Arteria_afectada|art. cerebral media
C0000017|_SUG_Arteria_afectada|ARTERIA VERTEBROBASILAR
C0000017|_SUG_Arteria_afectada|CEREBRALES POSTERIORES
C0000017|_SUG_Arteria_afectada|NO ESPECIF.
C0000017|_SUG_Arteria_afectada|vertebral
C0000002|_SUG_Ataque_isquemico_transitorio|AITs
C0000020|_SUG_Etiologia|cardioemebolico
C0000020|_SUG_Etiologia|CE
C0000020|_SUG_Etiologia|etiologia pendent de filiacio
C0000020|_SUG_Etiologia|hipertensivo
C0000020|_SUG_Etiologia|indeterminado (estudio incompleto)
C0000020|_SUG_Etiologia|insual
C0000020|_SUG_Etiologia|origen cardiaco
C0000019|_SUG_Lateralizacion|BIHEMISFERICO
C0000019|_SUG_Lateralizacion|dcho
C0000019|_SUG_Lateralizacion|derecho
C0000019|_SUG_Lateralizacion|ESQ.
C0000019|_SUG_Lateralizacion|IZDO
C0000018|_SUG_Localizacion|emporo-insular
C0000018|_SUG_Localizacion|fronto-occipital
C0000018|_SUG_Localizacion|frontal y occipital
C0000018|_SUG_Localizacion|gangliobasal
C0000018|_SUG_Localizacion|indeterminada
C0000018|_SUG_Localizacion|lenticulocapsular
C0000018|_SUG_Localizacion|lenticulocapsulotalamico
C0000018|_SUG_Localizacion|PROTUBERANCIAL
C0000018|_SUG_Localizacion|temporobasal
C0000018|_SUG_Localizacion|temporal basal
C0000018|_SUG_Localizacion|territorio indeterminado
C0000018|_SUG_Localizacion|ventricular
C0000021|_SUG_TAC_craneal|Tomografia axial computeritzada de cap
C0000007|_SUG_Test_de_disfagia|Test deglucion
C0000016|_SUG_Tratamiento_antiagregante|A.A.S.
C0000016|_SUG_Tratamiento_antiagregante|acetilsalicilico
C0000005|_SUG_Trombectomia_mecanica|terapia endovascular
C0000004|_SUG_Trombolisis_intravenosa|rTPA ev
C0000024|_SUG_Recanalizacion|Recanalizacion
C0000025|_SUG_Puerta_aguja|puerta aguja
