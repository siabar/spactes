c0000001|_SUG_Ictus_isquemico|Infarto
c0000001|_SUG_Ictus_isquemico|Avc
c0000001|_SUG_Ictus_isquemico|Avc isquemic
c0000001|_SUG_Ictus_isquemico|ICTUS ISQUÉMIC
c0000001|_SUG_Ictus_isquemico|ECVA isquémica
c0000001|_SUG_Ictus_isquemico|ECVA ISQUÉMICA
c0000001|_SUG_Ictus_isquemico|ECVA ISQUÉMICA: INFARTO
c0000001|_SUG_Ictus_isquemico|ECVA: INFARTOS ISQUÉMICOS
c0000001|_SUG_Ictus_isquemico|Ictus isquémico
c0000001|_SUG_Ictus_isquemico|Infart
c0000001|_SUG_Ictus_isquemico|Infart isquèmic
c0000001|_SUG_Ictus_isquemico|INFARTO
c0000001|_SUG_Ictus_isquemico|Infarto isquémico
c0000001|_SUG_Ictus_isquemico|Infarto isquémico
c0000001|_SUG_Ictus_isquemico|infarto isquémico
c0000001|_SUG_Ictus_isquemico|Infarto isquémico agudo
c0000001|_SUG_Ictus_isquemico|Infartos
c0000001|_SUG_Ictus_isquemico|Infartos isquémicos
c0000001|_SUG_Ictus_isquemico|sufusión hemorrágica
c0000001|_SUG_Ictus_isquemico|transformació hemorrágica
c0000001|_SUG_Ictus_isquemico|Transformacióhemorrágica
c0000001|_SUG_Ictus_isquemico|transformación hemorrágica
c0000002|_SUG_Ataque_isquemico_transitorio|ACCIDENTE TRANSITORI ISQUÉMICO.
c0000002|_SUG_Ataque_isquemico_transitorio|ictus
c0000002|_SUG_Ataque_isquemico_transitorio|ICTUS MINOR
c0000002|_SUG_Ataque_isquemico_transitorio|Infarto clínicamente regresivo
c0000002|_SUG_Ataque_isquemico_transitorio|Síndrome sensitivo-motor regresivo
c0000003|_SUG_Hemorragia_cerebral|AVC HEMORRAGIC
c0000003|_SUG_Hemorragia_cerebral|AVC HEMORRÀGIC
c0000003|_SUG_Hemorragia_cerebral|Hematoma
c0000003|_SUG_Hemorragia_cerebral|hematoma
c0000003|_SUG_Hemorragia_cerebral|HEMATOMA
c0000003|_SUG_Hemorragia_cerebral|Hemorragia
c0000003|_SUG_Hemorragia_cerebral|HEMORRAGIA
c0000003|_SUG_Hemorragia_cerebral|HEMORRAGIA PARENQUIMATOSA CEREBRAL MASIVA
c0000004|_SUG_Trombolisis_intravenosa|ECAS IV
c0000004|_SUG_Trombolisis_intravenosa|fibrinolítico
c0000004|_SUG_Trombolisis_intravenosa|fibrinolótico
c0000004|_SUG_Trombolisis_intravenosa|tPAev
c0000004|_SUG_Trombolisis_intravenosa|tractat amb firbinolisi
c0000004|_SUG_Trombolisis_intravenosa|tratamiento con alteplasa
c0000004|_SUG_Trombolisis_intravenosa|Tratamiento con RTPA
c0000004|_SUG_Trombolisis_intravenosa|tratamiento fibrinolítico
c0000004|_SUG_Trombolisis_intravenosa|trombolisis
c0000004|_SUG_Trombolisis_intravenosa|trombolisis
c0000005|_SUG_Trombectomia_mecanica|TEV
c0000005|_SUG_Trombectomia_mecanica|Trombectomíaendovascular
c0000005|_SUG_Trombectomia_mecanica|Trombectomiamecànica
c0000009|_SUG_NIHSS|NHISS 7
c0000009|_SUG_NIHSS|NIH 0
c0000009|_SUG_NIHSS|NIH 4
c0000009|_SUG_NIHSS|NIH 4)
c0000009|_SUG_NIHSS|NIH 8
c0000009|_SUG_NIHSS|NIH 9
c0000009|_SUG_NIHSS|NIH: 0
c0000009|_SUG_NIHSS|NIH: 0
c0000009|_SUG_NIHSS|NIH: 10
c0000009|_SUG_NIHSS|NIH: 7
c0000009|_SUG_NIHSS|NIH:1
c0000009|_SUG_NIHSS|NIH:12
c0000009|_SUG_NIHSS|NIH:16
c0000009|_SUG_NIHSS|NIH:3
c0000009|_SUG_NIHSS|NIH:3
c0000009|_SUG_NIHSS|NIH:6
c0000009|_SUG_NIHSS|NIH:8
c0000009|_SUG_NIHSS|NIHSS: 0-0-0-0- 0/0-0-0-0-0/0-0-0-1-0= 1
c0000009|_SUG_NIHSS|NIHSS=0
c0000009|_SUG_NIHSS|NIHSS=17
c0000009|_SUG_NIHSS|NIHSS=4
c0000009|_SUG_NIHSS|NISHSS=5
c0000009|_SUG_NIHSS|NISSH 14
c0000009|_SUG_NIHSS|PUNTUACION TOTAL NIH:19
c0000009|_SUG_NIHSS|PUNTUACION TOTAL NIH:6
c0000009|_SUG_NIHSS|NIHSS de 1
c0000010|_SUG_ASPECTS|ASPECTS 10
c0000010|_SUG_ASPECTS|ASPECTS (de 1 a 10): 10
c0000010|_SUG_ASPECTS|ASPECTS 6
c0000010|_SUG_ASPECTS|ASPECTS=10
c0000011|_SUG_mRankin|mRS 1-2
c0000011|_SUG_mRankin|mRS: 0
c0000011|_SUG_mRankin|MRS 0
c0000011|_SUG_mRankin|mRs:3
c0000011|_SUG_mRankin|mRs:3
c0000011|_SUG_mRankin|mRS=0
c0000011|_SUG_mRankin|mRs=0
c0000011|_SUG_mRankin|mRS=1
c0000011|_SUG_mRankin|mRS=1
c0000011|_SUG_mRankin|mRs=2
c0000011|_SUG_mRankin|mRS=2
c0000011|_SUG_mRankin|mRs=3
c0000011|_SUG_mRankin|mRS=3
c0000011|_SUG_mRankin|mRs=4
c0000011|_SUG_mRankin|mRS=4
c0000011|_SUG_mRankin|mRS=5
c0000011|_SUG_mRankin|mRs0
c0000011|_SUG_mRankin|mRS1
c0000011|_SUG_mRankin|mRS1
c0000011|_SUG_mRankin|mRS2
c0000011|_SUG_mRankin|mRS2
c0000011|_SUG_mRankin|Rankin:5
c0000011|_SUG_mRankin|Rankin=0
c0000011|_SUG_mRankin|Rankin0
c0000013|_SUG_Tratamiento_anticoagulante|Dabigatran
c0000015|_SUG_Tratamiento_antiagregante|AC ACETILSALICILICO
c0000015|_SUG_Tratamiento_antiagregante|Acido acetilsalicilico
c0000015|_SUG_Tratamiento_antiagregante|Acido acetilsalicílico
c0000015|_SUG_Tratamiento_antiagregante|Ácido acetilsalicílico
c0000015|_SUG_Tratamiento_antiagregante|ÁCIDO ACETILSALICÍLICO
c0000015|_SUG_Tratamiento_antiagregante|Ácido acetilsalicílico:
c0000015|_SUG_Tratamiento_antiagregante|Adiro
c0000015|_SUG_Tratamiento_antiagregante|Aspirina
c0000015|_SUG_Tratamiento_antiagregante|cido acetilsalicilico
c0000017|_SUG_Arteria_afectada|A.COROIDEA ANT
c0000017|_SUG_Arteria_afectada|A2
c0000017|_SUG_Arteria_afectada|ACA
c0000017|_SUG_Arteria_afectada|ACM
c0000017|_SUG_Arteria_afectada|art Vertebral
c0000017|_SUG_Arteria_afectada|arteria carotide
c0000017|_SUG_Arteria_afectada|arteria cerebral mitja
c0000017|_SUG_Arteria_afectada|artèria cerebral mitja
c0000017|_SUG_Arteria_afectada|ARTERIES CEREBRALS MITGES
c0000017|_SUG_Arteria_afectada|C1
c0000017|_SUG_Arteria_afectada|carótida primitiva
c0000017|_SUG_Arteria_afectada|carotidea
c0000017|_SUG_Arteria_afectada|CAROTÍDEA
c0000017|_SUG_Arteria_afectada|INDETERM I NA DO
c0000017|_SUG_Arteria_afectada|indeterminado
c0000017|_SUG_Arteria_afectada|M1-M2
c0000017|_SUG_Arteria_afectada|M2
c0000017|_SUG_Arteria_afectada|M3
c0000017|_SUG_Arteria_afectada|M4
c0000017|_SUG_Arteria_afectada|M5
c0000017|_SUG_Arteria_afectada|núcleo lenticular
c0000017|_SUG_Arteria_afectada|territorio indeterminado
c0000017|_SUG_Arteria_afectada|TICA
c0000017|_SUG_Arteria_afectada|V1
c0000017|_SUG_Arteria_afectada|VB
c0000017|_SUG_Arteria_afectada|VERTEBR BASILAR
c0000017|_SUG_Arteria_afectada|vertebro-basilar
c0000017|_SUG_Arteria_afectada|vertebrobasilar
c0000018|_SUG_Localizacion|BULBAR
c0000018|_SUG_Localizacion|càpsulo-talàmic
c0000018|_SUG_Localizacion|capsulotalamico
c0000018|_SUG_Localizacion|CAPSULOTALÁMICO
c0000018|_SUG_Localizacion|corona radiada
c0000018|_SUG_Localizacion|fronto-insular
c0000018|_SUG_Localizacion|fronto-temporo-insular
c0000018|_SUG_Localizacion|ganglicapsular
c0000018|_SUG_Localizacion|ganglios basales
c0000018|_SUG_Localizacion|GANGLIOS BASALES
c0000018|_SUG_Localizacion|INDETERM I NA DO
c0000018|_SUG_Localizacion|indeterminado
c0000018|_SUG_Localizacion|LACUNAR
c0000018|_SUG_Localizacion|lacunar
c0000018|_SUG_Localizacion|parcial
c0000018|_SUG_Localizacion|parietooccipital
c0000018|_SUG_Localizacion|profundes
c0000018|_SUG_Localizacion|subcorticals
c0000018|_SUG_Localizacion|talàmica
c0000018|_SUG_Localizacion|TALAMICO
c0000018|_SUG_Localizacion|talámico
c0000018|_SUG_Localizacion|talamo-capuslar
c0000018|_SUG_Localizacion|territorio indeterminado
c0000018|_SUG_Localizacion|ventriculos
c0000019|_SUG_Lateralizacion|ambas
c0000019|_SUG_Lateralizacion|bilateral
c0000019|_SUG_Lateralizacion|BILATERAL
c0000019|_SUG_Lateralizacion|bilaterales
c0000019|_SUG_Lateralizacion|BILATERALS
c0000019|_SUG_Lateralizacion|BILATERASL
c0000019|_SUG_Lateralizacion|D
c0000019|_SUG_Lateralizacion|derecha
c0000019|_SUG_Lateralizacion|DERECHOS
c0000019|_SUG_Lateralizacion|dret
c0000019|_SUG_Lateralizacion|dreta
c0000019|_SUG_Lateralizacion|DRETA
c0000019|_SUG_Lateralizacion|e
c0000019|_SUG_Lateralizacion|E
c0000019|_SUG_Lateralizacion|esq
c0000019|_SUG_Lateralizacion|esquerra
c0000019|_SUG_Lateralizacion|esquerre
c0000019|_SUG_Lateralizacion|esquerres
c0000019|_SUG_Lateralizacion|I
c0000019|_SUG_Lateralizacion|indeterminada
c0000019|_SUG_Lateralizacion|izda
c0000019|_SUG_Lateralizacion|IZQ
c0000019|_SUG_Lateralizacion|izquierda
c0000020|_SUG_Etiologia|a estudio
c0000020|_SUG_Etiologia|ateromatosis
c0000020|_SUG_Etiologia|Cavernoma de circunvolución
c0000020|_SUG_Etiologia|Criptogènic
c0000020|_SUG_Etiologia|criptogénico
c0000020|_SUG_Etiologia|Disecció
c0000020|_SUG_Etiologia|embòlic
c0000020|_SUG_Etiologia|embólico
c0000020|_SUG_Etiologia|embólico
c0000020|_SUG_Etiologia|indeterminada (posiblemente paraneoplásico)
c0000020|_SUG_Etiologia|infrecuente
c0000020|_SUG_Etiologia|LACUNAR
c0000020|_SUG_Etiologia|lacunar
c0000020|_SUG_Etiologia|malformación arteriovenosa
c0000020|_SUG_Etiologia|mecanisme embòlic
c0000021|_SUG_TAC_craneal|AgioTAC
c0000021|_SUG_TAC_craneal|TA C crani al
c0000021|_SUG_TAC_craneal|TAC
c0000021|_SUG_TAC_craneal|TAC cerebral
c0000021|_SUG_TAC_craneal|Tac de cráneo
c0000021|_SUG_TAC_craneal|TC
c0000021|_SUG_TAC_craneal|Tc craneal
c0000021|_SUG_TAC_craneal|Tc cranial