C0000001|_SUG_Ictus_isquemico|ictus isquémico
C0000001|_SUG_Ictus_isquemico|ictus
C0000001|_SUG_Ictus_isquemico|infarto cerebral
C0000001|_SUG_Ictus_isquemico|accidente cerebrovascular
C0000001|_SUG_Ictus_isquemico|ictus isquémico con transformación hemorrágica
C0000001|_SUG_Ictus_isquemico|AVC
C0000002|_SUG_Ataque_isquemico_transitorio|ataque isquémico transitorio
C0000002|_SUG_Ataque_isquemico_transitorio|AIT
C0000002|_SUG_Ataque_isquemico_transitorio|TIA
C0000003|_SUG_Hemorragia_cerebral|hemorragia cerebral
C0000003|_SUG_Hemorragia_cerebral|hemorragia intracerebral
C0000003|_SUG_Hemorragia_cerebral|ictus hemorrágico
C0000003|_SUG_Hemorragia_cerebral|hematoma cerebral
C0000004|_SUG_Trombolisis_intravenosa|trombólisis intravenosa
C0000004|_SUG_Trombolisis_intravenosa|fibrinolisis
C0000004|_SUG_Trombolisis_intravenosa|rtPA
C0000004|_SUG_Trombolisis_intravenosa|fibrinolisis iv
C0000004|_SUG_Trombolisis_intravenosa|fibrinolisis endovenosa
C0000004|_SUG_Trombolisis_intravenosa|tratamiento trombolítico
C0000004|_SUG_Trombolisis_intravenosa|fibrinólisis sistémica con rtPA ev
C0000005|_SUG_Trombectomia_mecanica|tratamiento endovascular
C0000005|_SUG_Trombectomia_mecanica|trombectomía
C0000005|_SUG_Trombectomia_mecanica|trombectomía mecánica
C0000006|_SUG_Trombolisis_intraarterial|trombólisis ia
C0000006|_SUG_Trombolisis_intraarterial|trombólisis intraarterial
C0000007|_SUG_Test_de_disfagia|test de disfagia
C0000007|_SUG_Test_de_disfagia|test de deglución
C0000008|_SUG_mRankin_previa|Escala de Rankin modificada 0
C0000008|_SUG_mRankin_previa|mRankin 0
C0000008|_SUG_mRankin_previa|Rankin 0
C0000008|_SUG_mRankin_previa|mRs 0
C0000008|_SUG_mRankin_previa|mRS 0
C0000009|_SUG_NIHSS_previa|Escala NIHSS 0
C0000009|_SUG_NIHSS_previa|NIHSS 0
C0000010|_SUG_ASPECTS|escala ASPECTS 0
C0000010|_SUG_ASPECTS|ASPECTS score 0
C0000010|_SUG_ASPECTS|ASPECTS 0
C0000011|_SUG_mRankin_alta|Escala de Rankin modificada 0
C0000011|_SUG_mRankin_alta|mRankin 0
C0000011|_SUG_mRankin_alta|Rankin 0
C0000011|_SUG_mRankin_alta|mRS 0
C0000011|_SUG_mRankin_alta|mRs 0
C0000012|_SUG_NIHSS_alta|Escala NIHSS 0
C0000012|_SUG_NIHSS_alta|NIHSS 0
C0000013|_SUG_Tratamiento_anticoagulante_hab|acenocumarol
C0000013|_SUG_Tratamiento_anticoagulante_hab|warfarin
C0000013|_SUG_Tratamiento_anticoagulante_hab|heparin
C0000013|_SUG_Tratamiento_anticoagulante_hab|dalteparin
C0000013|_SUG_Tratamiento_anticoagulante_hab|enoxaparin
C0000013|_SUG_Tratamiento_anticoagulante_hab|nadroparin
C0000013|_SUG_Tratamiento_anticoagulante_hab|parnaparin
C0000013|_SUG_Tratamiento_anticoagulante_hab|reviparin
C0000013|_SUG_Tratamiento_anticoagulante_hab|bemiparin
C0000013|_SUG_Tratamiento_anticoagulante_hab|dabigatran etexilate
C0000013|_SUG_Tratamiento_anticoagulante_hab|rivaroxaban
C0000013|_SUG_Tratamiento_anticoagulante_hab|apixaban
C0000013|_SUG_Tratamiento_anticoagulante_hab|edoxaban
C0000013|_SUG_Tratamiento_anticoagulante_hab|B01AA07
C0000013|_SUG_Tratamiento_anticoagulante_hab|B01AA03
C0000013|_SUG_Tratamiento_anticoagulante_hab|B01AB01
C0000013|_SUG_Tratamiento_anticoagulante_hab|B01AB04
C0000013|_SUG_Tratamiento_anticoagulante_hab|B01AB05
C0000013|_SUG_Tratamiento_anticoagulante_hab|B01AB06
C0000013|_SUG_Tratamiento_anticoagulante_hab|B01AB07
C0000013|_SUG_Tratamiento_anticoagulante_hab|B01AB08
C0000013|_SUG_Tratamiento_anticoagulante_hab|B01AB12
C0000013|_SUG_Tratamiento_anticoagulante_hab|B01AE07
C0000013|_SUG_Tratamiento_anticoagulante_hab|B01AF01
C0000013|_SUG_Tratamiento_anticoagulante_hab|B01AF02
C0000013|_SUG_Tratamiento_anticoagulante_hab|B01AF03
C0000013|_SUG_Tratamiento_anticoagulante_hab|sintrom
C0000013|_SUG_Tratamiento_anticoagulante_hab|aldocumar
C0000013|_SUG_Tratamiento_anticoagulante_hab|Heparina
C0000013|_SUG_Tratamiento_anticoagulante_hab|fragmin
C0000013|_SUG_Tratamiento_anticoagulante_hab|clexane
C0000013|_SUG_Tratamiento_anticoagulante_hab|fraxiparina
C0000013|_SUG_Tratamiento_anticoagulante_hab|hibor
C0000013|_SUG_Tratamiento_anticoagulante_hab|pradaxa
C0000013|_SUG_Tratamiento_anticoagulante_hab|xarelto
C0000013|_SUG_Tratamiento_anticoagulante_hab|eliquis
C0000013|_SUG_Tratamiento_anticoagulante_hab|lixiana
C0000014|_SUG_Tratamiento_anticoagulante_alta|acenocumarol
C0000014|_SUG_Tratamiento_anticoagulante_alta|warfarin
C0000014|_SUG_Tratamiento_anticoagulante_alta|heparin
C0000014|_SUG_Tratamiento_anticoagulante_alta|dalteparin
C0000014|_SUG_Tratamiento_anticoagulante_alta|enoxaparin
C0000014|_SUG_Tratamiento_anticoagulante_alta|nadroparin
C0000014|_SUG_Tratamiento_anticoagulante_alta|parnaparin
C0000014|_SUG_Tratamiento_anticoagulante_alta|reviparin
C0000014|_SUG_Tratamiento_anticoagulante_alta|bemiparin
C0000014|_SUG_Tratamiento_anticoagulante_alta|dabigatran etexilate
C0000014|_SUG_Tratamiento_anticoagulante_alta|rivaroxaban
C0000014|_SUG_Tratamiento_anticoagulante_alta|apixaban
C0000014|_SUG_Tratamiento_anticoagulante_alta|edoxaban
C0000014|_SUG_Tratamiento_anticoagulante_alta|B01AA07
C0000014|_SUG_Tratamiento_anticoagulante_alta|B01AA03
C0000014|_SUG_Tratamiento_anticoagulante_alta|B01AB01
C0000014|_SUG_Tratamiento_anticoagulante_alta|B01AB04
C0000014|_SUG_Tratamiento_anticoagulante_alta|B01AB05
C0000014|_SUG_Tratamiento_anticoagulante_alta|B01AB06
C0000014|_SUG_Tratamiento_anticoagulante_alta|B01AB07
C0000014|_SUG_Tratamiento_anticoagulante_alta|B01AB08
C0000014|_SUG_Tratamiento_anticoagulante_alta|B01AB12
C0000014|_SUG_Tratamiento_anticoagulante_alta|B01AE07
C0000014|_SUG_Tratamiento_anticoagulante_alta|B01AF01
C0000014|_SUG_Tratamiento_anticoagulante_alta|B01AF02
C0000014|_SUG_Tratamiento_anticoagulante_alta|B01AF03
C0000014|_SUG_Tratamiento_anticoagulante_alta|sintrom
C0000014|_SUG_Tratamiento_anticoagulante_alta|aldocumar
C0000014|_SUG_Tratamiento_anticoagulante_alta|Heparina
C0000014|_SUG_Tratamiento_anticoagulante_alta|fragmin
C0000014|_SUG_Tratamiento_anticoagulante_alta|clexane
C0000014|_SUG_Tratamiento_anticoagulante_alta|fraxiparina
C0000014|_SUG_Tratamiento_anticoagulante_alta|hibor
C0000014|_SUG_Tratamiento_anticoagulante_alta|pradaxa
C0000014|_SUG_Tratamiento_anticoagulante_alta|xarelto
C0000014|_SUG_Tratamiento_anticoagulante_alta|eliquis
C0000014|_SUG_Tratamiento_anticoagulante_alta|lixiana
C0000015|_SUG_Tratamiento_antiagregante_hab|clopidogrel
C0000015|_SUG_Tratamiento_antiagregante_hab|ticlopidine
C0000015|_SUG_Tratamiento_antiagregante_hab|acetylsalicylic acid
C0000015|_SUG_Tratamiento_antiagregante_hab|dipyridamole
C0000015|_SUG_Tratamiento_antiagregante_hab|abciximab
C0000015|_SUG_Tratamiento_antiagregante_hab|tirofiban
C0000015|_SUG_Tratamiento_antiagregante_hab|triflusal
C0000015|_SUG_Tratamiento_antiagregante_hab|cilostazol
C0000015|_SUG_Tratamiento_antiagregante_hab|ticagrelor
C0000015|_SUG_Tratamiento_antiagregante_hab|cangrelor
C0000015|_SUG_Tratamiento_antiagregante_hab|prasugler
C0000015|_SUG_Tratamiento_antiagregante_hab|combinations
C0000015|_SUG_Tratamiento_antiagregante_hab|acetylsalicylic acid, combinations with proton pump inhibitors
C0000015|_SUG_Tratamiento_antiagregante_hab|B01AC04
C0000015|_SUG_Tratamiento_antiagregante_hab|B01AC05
C0000015|_SUG_Tratamiento_antiagregante_hab|B01AC06
C0000015|_SUG_Tratamiento_antiagregante_hab|B01AC07
C0000015|_SUG_Tratamiento_antiagregante_hab|B01AC13
C0000015|_SUG_Tratamiento_antiagregante_hab|B01AC17
C0000015|_SUG_Tratamiento_antiagregante_hab|B01AC18
C0000015|_SUG_Tratamiento_antiagregante_hab|B01AC23
C0000015|_SUG_Tratamiento_antiagregante_hab|B01AC24
C0000015|_SUG_Tratamiento_antiagregante_hab|B01AC25
C0000015|_SUG_Tratamiento_antiagregante_hab|B01AC22
C0000015|_SUG_Tratamiento_antiagregante_hab|B01AC30
C0000015|_SUG_Tratamiento_antiagregante_hab|B01AC56
C0000015|_SUG_Tratamiento_antiagregante_hab|plavix
C0000015|_SUG_Tratamiento_antiagregante_hab|tiklid
C0000015|_SUG_Tratamiento_antiagregante_hab|Adiro
C0000015|_SUG_Tratamiento_antiagregante_hab|AAS
C0000015|_SUG_Tratamiento_antiagregante_hab|persantin
C0000015|_SUG_Tratamiento_antiagregante_hab|reopro
C0000015|_SUG_Tratamiento_antiagregante_hab|agrastat
C0000015|_SUG_Tratamiento_antiagregante_hab|disgren
C0000015|_SUG_Tratamiento_antiagregante_hab|ekistol
C0000015|_SUG_Tratamiento_antiagregante_hab|pletal
C0000015|_SUG_Tratamiento_antiagregante_hab|brilique
C0000016|_SUG_Tratamiento_antiagregante_alta|clopidogrel
C0000016|_SUG_Tratamiento_antiagregante_alta|ticlopidine
C0000016|_SUG_Tratamiento_antiagregante_alta|acetylsalicylic acid
C0000016|_SUG_Tratamiento_antiagregante_alta|dipyridamole
C0000016|_SUG_Tratamiento_antiagregante_alta|abciximab
C0000016|_SUG_Tratamiento_antiagregante_alta|tirofiban
C0000016|_SUG_Tratamiento_antiagregante_alta|triflusal
C0000016|_SUG_Tratamiento_antiagregante_alta|cilostazol
C0000016|_SUG_Tratamiento_antiagregante_alta|ticagrelor
C0000016|_SUG_Tratamiento_antiagregante_alta|cangrelor
C0000016|_SUG_Tratamiento_antiagregante_alta|prasugler
C0000016|_SUG_Tratamiento_antiagregante_alta|combinations
C0000016|_SUG_Tratamiento_antiagregante_alta|acetylsalicylic acid, combinations with proton pump inhibitors
C0000016|_SUG_Tratamiento_antiagregante_alta|B01AC04
C0000016|_SUG_Tratamiento_antiagregante_alta|B01AC05
C0000016|_SUG_Tratamiento_antiagregante_alta|B01AC06
C0000016|_SUG_Tratamiento_antiagregante_alta|B01AC07
C0000016|_SUG_Tratamiento_antiagregante_alta|B01AC13
C0000016|_SUG_Tratamiento_antiagregante_alta|B01AC17
C0000016|_SUG_Tratamiento_antiagregante_alta|B01AC18
C0000016|_SUG_Tratamiento_antiagregante_alta|B01AC23
C0000016|_SUG_Tratamiento_antiagregante_alta|B01AC24
C0000016|_SUG_Tratamiento_antiagregante_alta|B01AC25
C0000016|_SUG_Tratamiento_antiagregante_alta|B01AC22
C0000016|_SUG_Tratamiento_antiagregante_alta|B01AC30
C0000016|_SUG_Tratamiento_antiagregante_alta|B01AC56
C0000016|_SUG_Tratamiento_antiagregante_alta|plavix
C0000016|_SUG_Tratamiento_antiagregante_alta|tiklid
C0000016|_SUG_Tratamiento_antiagregante_alta|Adiro
C0000016|_SUG_Tratamiento_antiagregante_alta|AAS
C0000016|_SUG_Tratamiento_antiagregante_alta|persantin
C0000016|_SUG_Tratamiento_antiagregante_alta|reopro
C0000016|_SUG_Tratamiento_antiagregante_alta|agrastat
C0000016|_SUG_Tratamiento_antiagregante_alta|disgren
C0000016|_SUG_Tratamiento_antiagregante_alta|ekistol
C0000016|_SUG_Tratamiento_antiagregante_alta|pletal
C0000016|_SUG_Tratamiento_antiagregante_alta|brilique
C0000017|_SUG_Arteria_afectada|Arteria carótida común
C0000017|_SUG_Arteria_afectada|ACC
C0000017|_SUG_Arteria_afectada|Arteria carótida interna
C0000017|_SUG_Arteria_afectada|ACI
C0000017|_SUG_Arteria_afectada|Arteria carótida interna terminal
C0000017|_SUG_Arteria_afectada|ACI-T
C0000017|_SUG_Arteria_afectada|AICA
C0000017|_SUG_Arteria_afectada|Arteria cerebral media
C0000017|_SUG_Arteria_afectada|ACM
C0000017|_SUG_Arteria_afectada|Arteria cerebral media segmento M1
C0000017|_SUG_Arteria_afectada|M1
C0000017|_SUG_Arteria_afectada|Arteria cerebral media segmento M2
C0000017|_SUG_Arteria_afectada|M2
C0000017|_SUG_Arteria_afectada|Arteria cerebral anterior
C0000017|_SUG_Arteria_afectada|ACA
C0000017|_SUG_Arteria_afectada|Arteria cerebral posterior
C0000017|_SUG_Arteria_afectada|ACP
C0000017|_SUG_Arteria_afectada|Arteria lenticuloestriada
C0000017|_SUG_Arteria_afectada|Arteria coroidea anterior
C0000017|_SUG_Arteria_afectada|Arteria coroidea posterior
C0000017|_SUG_Arteria_afectada|Arteria cerebelosa superior
C0000017|_SUG_Arteria_afectada|ACS
C0000017|_SUG_Arteria_afectada|Arteria cerebelosa anteroinferior
C0000017|_SUG_Arteria_afectada|AICA
C0000017|_SUG_Arteria_afectada|Arteria cerebelosa posteroinferior
C0000017|_SUG_Arteria_afectada|PICA
C0000017|_SUG_Arteria_afectada|Arteria vertebral
C0000017|_SUG_Arteria_afectada|Arteria basilar
C0000017|_SUG_Arteria_afectada|AB
C0000018|_SUG_Localizacion|Infarto total de circulación anterior
C0000018|_SUG_Localizacion|TACI
C0000018|_SUG_Localizacion|Infarto parcial de circulación anterior
C0000018|_SUG_Localizacion|PACI
C0000018|_SUG_Localizacion|Infarto lacunar
C0000018|_SUG_Localizacion|LACI
C0000018|_SUG_Localizacion|Infarto de circulación posterior
C0000018|_SUG_Localizacion|POCI
C0000018|_SUG_Localizacion|Lobar
C0000018|_SUG_Localizacion|frontal 
C0000018|_SUG_Localizacion|cortical
C0000018|_SUG_Localizacion|temporal 
C0000018|_SUG_Localizacion|parietal 
C0000018|_SUG_Localizacion|occipital
C0000018|_SUG_Localizacion|profunda 
C0000018|_SUG_Localizacion|ggbb
C0000018|_SUG_Localizacion|ganglios de la base
C0000018|_SUG_Localizacion|tálamo 
C0000018|_SUG_Localizacion|putamen 
C0000018|_SUG_Localizacion|caudado 
C0000018|_SUG_Localizacion|lenticular 
C0000018|_SUG_Localizacion|pálido
C0000018|_SUG_Localizacion|Intraventricular
C0000018|_SUG_Localizacion|posterior
C0000018|_SUG_Localizacion|tronco
C0000018|_SUG_Localizacion|cerebelosa
C0000019|_SUG_Lateralizacion|Izquierda
C0000019|_SUG_Lateralizacion|Izq
C0000019|_SUG_Lateralizacion|I
C0000019|_SUG_Lateralizacion|Derecha
C0000019|_SUG_Lateralizacion|Dcha
C0000019|_SUG_Lateralizacion|D
C0000019|_SUG_Lateralizacion|Tronco cerebral 
C0000020|_SUG_Etiologia|Aterotrombótico
C0000020|_SUG_Etiologia|aterosclerótico
C0000020|_SUG_Etiologia|Cardioembólico
C0000020|_SUG_Etiologia|Lacunar
C0000020|_SUG_Etiologia|Indeterminado
C0000020|_SUG_Etiologia|ESUS
C0000020|_SUG_Etiologia|Indeterminado de causa doble
C0000020|_SUG_Etiologia|Indeterminado por estudio incompleto
C0000020|_SUG_Etiologia|Inhabitual
C0000020|_SUG_Etiologia|Hipertensiva
C0000020|_SUG_Etiologia|angiopatía amiloide
C0000020|_SUG_Etiologia|secundaria a malformación vascular
C0000020|_SUG_Etiologia|aneurisma
C0000020|_SUG_Etiologia|secundaria a tumor
C0000020|_SUG_Etiologia|indeterminada
C0000021|_SUG_TAC_craneal|TAC craneal
C0000021|_SUG_TAC_craneal|TC craneal
C0000021|_SUG_TAC_craneal|TC cranial
C0000021|_SUG_TAC_craneal|TC de cráneo
C0000021|_SUG_TAC_craneal|TC